library ieee;
use ieee.std_logic_1164.all;

entity Register_Module is
port(
	